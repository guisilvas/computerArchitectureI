// CI - Standard logic
// Full-Custom IC (uses transistor)
//FPGA

// Gates : AND, OR, XOR, NOT
// Muxes/Demuxes
// Registers/Memory
// Aithmetic Operations (Adder, Sbtracter, Multiplier, etc)
// State Machines
// Any combinations of Above

module

end module
